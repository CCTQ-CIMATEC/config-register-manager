package bus_definitions;

localparam DATA_WIDTH = 32;
localparam ADDR_WIDTH = 32;

endpackage: bus_definitions